module ttt (
    input  a,
    output b
);
//심심해
endmodule
