module ttt (
    input  a,
    output b
);
endmodule
